`include "agent1_config.sv"
`include "agent2_config.sv"
`include "env_config.sv"

`include "xtn1.sv"
`include "xtn2.sv"

`include "driver1.sv"
`include "monitor1.sv"
`include "agent1.sv"

`include "driver2.sv"
`include "monitor2.sv"
`include "agent2.sv"

`include "environment.sv"
`include "test.sv"